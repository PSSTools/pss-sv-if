
package psv_dpi;
    import psv::*;
endpackage

package pss_sv_if;

endpackage
